module priority_encoder;
endmodule
